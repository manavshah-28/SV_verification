interface intf(input logic clk);
 logic Stream;
 logic Tone;
 logic [2:0]Count;
endinterface 